module JK_FF(input J, K, Clk, R, En, output reg Q, output Qn);



endmodule //JK_FF

module JK_FF_tb();








endmodule //testbench